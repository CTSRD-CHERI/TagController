/* Copyright 2015 Matthew Naylor
 * All rights reserved.
 *
 * This software was developed by SRI International and the University of
 * Cambridge Computer Laboratory under DARPA/AFRL contract FA8750-10-C-0237
 * ("CTSRD"), as part of the DARPA CRASH research programme.
 *
 * This software was developed by SRI International and the University of
 * Cambridge Computer Laboratory under DARPA/AFRL contract FA8750-11-C-0249
 * ("MRC2"), as part of the DARPA MRC research programme.
 *
 * This software was developed by the University of Cambridge Computer
 * Laboratory as part of the Rigorous Engineering of Mainstream
 * Systems (REMS) project, funded by EPSRC grant EP/K008528/1.
 * 
 * This software was developed by SRI International and the University of
 * Cambridge Computer Laboratory (Department of Computer Science and
 * Technology) under DARPA contract HR0011-18-C-0016 ("ECATS"), as part of the
 * DARPA SSITH research programme.
 *
 * @BERI_LICENSE_HEADER_START@
 *
 * Licensed to BERI Open Systems C.I.C. (BERI) under one or more contributor
 * license agreements.  See the NOTICE file distributed with this work for
 * additional information regarding copyright ownership.  BERI licenses this
 * file to you under the BERI Hardware-Software License, Version 1.0 (the
 * "License"); you may not use this file except in compliance with the
 * License.  You may obtain a copy of the License at:
 *
 *   http://www.beri-open-systems.org/legal/license-1-0.txt
 *
 * Unless required by applicable law or agreed to in writing, Work distributed
 * under the License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
 * CONDITIONS OF ANY KIND, either express or implied.  See the License for the
 * specific language governing permissions and limitations under the License.
 *
 * @BERI_LICENSE_HEADER_END@
 */

import MemoryClient :: *;
import Vector       :: *;
import BlueCheck    :: *;
import StmtFSM      :: *;
import Memory       :: *;
import Clocks       :: *;
import FIFOF        :: *;
import Assert       :: *;
import Printf       :: *;

// ============================================================================
// Single-core
// ============================================================================

// Test equivalance against the golden model.
module [BlueCheck] checkSingle#( MemoryClient core
                               , MemoryClient gold
                               ) ();

  Reg#(Bool) init <- mkReg(True);
  
  let ensure <- mkEnsure;
  
  function Action setSameAddrMap(AddrMap map) =
    action
      core.setAddrMap(map);
      gold.setAddrMap(map);
    endaction;

  pre("setAddrMap", setSameAddrMap);
  equivf(3, "load" , core.load , gold.load);
  equivf(3, "store", core.store, gold.store);
  equivf(3, "getResponse", core.getResponse, gold.getResponse);

  // Read command-line arguments
  rule initialise (init);
    init <= False;
  endrule

endmodule
